* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)
*
* Experiment c. 3:
* pulzni odezva
*
* NOTES:
* - uzel 'in' byl prejmenovan na '3', z duvodu chyby .noise

*** NETLIST ***
Vin     3   0    5    PULSE 0 5 1u 1f 1f 5u 10u
Rb      a3  kat 1k
Rload 3   col {valrload}  ;stejne jako exp. 1a
Rs ref 0   100  ;Iout = Vref / Rs -> Rs = 32.5/10m
Xref    ref  0   kat TL431
Q1      col kat ref Q2N2222

Vrb     3   a3   0

*** PRIKAZY ***
.param valrload = 100 
.tran 8n 8u 0 10u SKIPBP
.lib tl431.mod
.lib MPS.lib
.probe
.op
.end
