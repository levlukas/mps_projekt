Zdroj proudu s vhodnou napetovou referenci

*** NETLIST ***
Vcc out 1 5  ;prozatim 5V
Rb out 4 100  ;prozatimni hodnota
Rload out 2 100  ;prozatimni hodnota
Rs 3 0 100  ;prozatimni hodnota
Xref 3 0 4 TL431  ;referenci napeti podle nahradniho obvodu
Q1 3 4 2 Q2N2222  ;nahodny jfet

Vaux 2 5 0  ; pomocne napeti pro vystup

*** PRIKAZY ***
.include /home/llev/OneDrive/4_letni/MPS/mps_projekt/tl431.mod
.lib mps.lib
.tran 10u 10m
.end
