* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)
*
* Experiment è. 2:
* Analyzujte spektrální hustotu umového výkonu a proudu zátìí
* v kmitoètovém pásmu 1 Hz a 150 kHz. Zjistìte efektivní hodnotu
* umového proudu v tomto frekvenèním pásmu (a srovnejte ji
* s velikostí pracovního proudu Iout).
*
* NOTES:
* - uzel 'in' byl prejmenovan na '3', z duvodu chyby .noise

*** NETLIST ***
Vin 3 0 1V  AC 5V  ;pro op 1V pro ac 5V bez phi0
Rb 3 kat 1k
Rload 3 col 100  ;stejne jako exp. 1a
Rs ref 0 100  ;Iout = Vref / Rs -> Rs = 2.5/25m
Xref ref 0 kat TL431
Q1 col kat ref Q2N2222


*** PRIKAZY ***
.lib ../tl431.mod
.lib ../MPS.lib
*.ac dec 1000 1 150k  ;ac analyza pro tisic bodu v def. freq
.noise V(3,col) Vin dec 1000 1 150k  ;pro LTspice bez AC
*.probe
.end
