* Experiment č. 1:
* Změřte teplotní koeficient proudu Iout při zátěži 100 Ω
* a Vcc = 5 V. Zjistěte závislost proudu Iout na velikosti
* zátěže. Ověřte výpočtem maximální hodnotu zátěže, kterou
* ještě může protékat nastavený konstantní proud.
*
* Experiment 1a:
* Změřte teplotní koeficient proudu Iout při zátěži 100 Ω
* a Vcc = 5 V.

*** NETLIST ***
Vcc out 0 5  ;prozatim 5V
Rb out 4 100  ;prozatimni hodnota
Rload out 2 100  ;prozatimni hodnota
Rs 3 0 100  ;prozatimni hodnota
Xref 3 0 4 TL431  ;referenci napeti podle nahradniho obvodu
Q1 3 4 2 Q2N2222

Vaux 2 5 0  ; pomocne napeti pro vystup

*** PRIKAZY ***
.include tl431.mod
.include mps.lib
.op
.end

