* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)
*
* Experiment c. 3:
* Sledovani ustalovani
*
* NOTES:
* - uzel 'in' byl prejmenovan na '3', z duvodu chyby .noise

*** NETLIST ***
*Vin 3 0 SIN 0 1 1k 0 0 0
Vin 3 0 PULSE 0 1 0 1f 1f {t0} {2*t0}
Rb 3 kat 1k
Rload 3 col 100  ;stejne jako exp. 1a
Rs ref 0 100  ;Iout = Vref / Rs -> Rs = 2.5/25m
Xref ref 0 kat TL431
Q1 col kat ref Q2N2222

*** PRIKAZY ***
.param t0=3u
.lib tl431.mod
.lib MPS.lib
.tran 1n 6u 0 0.1n SKIPBP
.probe  V(3) V(3,col) I(Rload)
.op
.end
