* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)
*
* Experiment č. 2:
* Analyzujte spektrální hustotu šumového výkonu a proudu
* zátěží v kmitočtovém pásmu 1 Hz až 150 kHz. Zjistěte
* efektivní hodnotu šumového proudu v tomto frekvenčním
* pásmu (a srovnejte ji s velikostí pracovního proudu Iout).


*** NETLIST ***
Vcc in 0 1V  AC 5V 0deg; pro op 1V, pro ac 5V bez phi0
Rb in kat 1k
Rload in col 100  ;stejne jako exp. 1a
Rs ref 0 100  ;Iout = Vref / Rs -> Rs = 2.5/25m
Xref ref 0 kat TL431
Q1 col kat ref Q2N2222


*** PRIKAZY ***
.include ../tl431.mod
.include ../MPS.lib
.op
*.ac dec 1000 1 150k  ;ac analyza pro tisic bodu v def. freq
.noise V(in,col) VCC dec 1000 1 150k
.end
