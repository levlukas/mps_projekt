* Experiment č. 1:
* Změřte teplotní koeficient proudu Iout při zátěži 100 Ω
* a Vcc = 5 V. Zjistěte závislost proudu Iout na velikosti
* zátěže. Ověřte výpočtem maximální hodnotu zátěže, kterou
* ještě může protékat nastavený konstantní proud.
*
* Experiment 1a:
* Změřte teplotní koeficient proudu Iout při zátěži 100 Ω
* a Vcc = 5 V.

*** NETLIST ***
Vcc in 0 sine(0 5 1k)  ;prozatim 5V
Rb auxib 4 15k  ;aby Ib=.25mA
Rload in 2 100  ;prozatimni hodnota
Rs 3 0 100  ;prozatimni hodnota
Xref 3 0 4 TL431  ;referenci napeti podle nahradniho obvodu
Q1 3 4 2 Q2N2222

Vaux 2 5 0  ; pomocne napeti pro vystup
VIb in auxib 0  ;pomocne pro Ib

*** PRIKAZY ***
.include tl431.mod
.op
.include MPS.lib
.tran 2u 2m
.end

