* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)

*** NETLIST ***
Vcc in 0 sine(0 5 1k)  ;prozatim 5Vpp
Rb auxib kat 15k  ;aby Ib=~250uA
Rload in col 100
Rs ref 0 100  ;prozatimni hodnota
Xref ref 0 kat TL431  ;referenci napeti podle nahradniho obvodu
Q1 col kat ref Q2N2222

VIb in auxib 0  ;pomocne pro Ib

*** PRIKAZY ***
.include tl431.mod
.op
.include MPS.lib
.tran 2u 2m
.end
