* ====== Zdroj proudu s vhodnou napetovou referenci ======
*
* Zvoleno: Iout = 25 mA
* Iout = Vref / Rs
* Rb = (Vcc - Vref - Vbe) / (Iout/h_fe + I_u1)
*
* Experiment č. 1:
* Změřte teplotní koeficient proudu Iout při zátěži 100 Ω a
* Vcc = 5 V. Zjistěte závislost proudu Iout na velikosti zátěže.
* Ověřte výpočtem maximální hodnotu zátěže, kterou ještě
* může protékat nastavený konstantní proud.
*
* Experiment 1b:
* Zjistěte závislost proudu Iout na velikosti zátěže.


*** NETLIST ***
Vcc 		in 		0 		{vccval}
Rb 		auxib 	kat	1k
Rload auxcol col 	{valRload}
Rs 		ref 		0 		100  ;Iout = Vref / Rs -> Rs = 2.5/25m
Xref 	ref 		0 		auxkat 	TL431
Q1 		col 		kat 	ref 			Q2N2222

* pomocne zdroje pro odecet proudu
VIb		in 	auxib 		0
Vka 	kat 	auxkat 	0
Vload 	in		auxcol		0


*** PRIKAZY ***
.op
.step param valrload 5 10k 100
.step param vccval list 5 15 36
.lib ../tl431.mod
.lib ../MPS.lib
.end
